module test (
    ports
);
    
endmodule